library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sumador is

port( 
	A: in std_logic_ ;
	B: in std_logic ;
	S: out std_logic ;
	Cs: out std_logic  );

end;

architecture behavioral of sumador is
begin

end behavioral;

